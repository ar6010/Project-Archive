--Andrew Ramirez

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;


entity adder is
port(
	A: in std_logic_vector(31 downto 0);
	B: in std_logic_vector(31 downto 0);
	S: out std_logic_vector(31 downto 0)
);
end entity adder;

architecture df of adder is

begin

	S <= A+B;

end architecture df;